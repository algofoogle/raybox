// SPDX-FileCopyrightText: 2023 Anton Maurovic <anton@maurovic.com>
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0


`default_nettype none
`timescale 1ns / 1ps

module trace_buffer(
    input       clk,
    input       cs,
    input       we,
    input       oe,
    input [9:0] column,

    inout [7:0] height, //SMELL: Should we have separate read/write ports for simplicity?
    inout       side
);

    reg [7:0]   height_out;
    reg         side_out;

    reg [7:0]   dummy_memory [0:640*2-1];
    initial $readmemh("assets/traces_capture_0001.hex", dummy_memory);

    // Tri-state buffer control for output mode:
    wire read_mode = (cs && oe && !we);
    assign height   = read_mode ? height_out    : 8'bz;
    assign side     = read_mode ? side_out      : 1'bz;

    // Memory write block:
    // ...TBC!...

    // Memory read block:
    always @(posedge clk) begin : MEM_READ
        if (read_mode) begin
            height_out = dummy_memory[{column,1'b0}];
            side_out = dummy_memory[{column,1'b1}][0];
        end
    end

endmodule
