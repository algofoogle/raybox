// Leading Zeroes Counter logic, borrowed from:
// https://github.com/ameetgohil/leading-zeroes-counter/blob/master/rtl/lzc.sv
// ...then fudged to just be Verilog (instead of SystemVerilog) and work with 32-bit input only.


module lzc #(
    parameter WIDTH=32 //SMELL: Not used.
)(
    input   [15:-16]    i_data,
    output   [5:0]      lzc_cnt
);

    function [5:0] f_lzc(input [15:-16] data);
        casez(data)
            32'b0:                                  f_lzc = 32;
            32'b1:                                  f_lzc = 31;
            32'b1?:                                 f_lzc = 30;
            32'b1??:                                f_lzc = 29;
            32'b1???:                               f_lzc = 28;
            32'b1????:                              f_lzc = 27;
            32'b1?????:                             f_lzc = 26;
            32'b1??????:                            f_lzc = 25;
            32'b1???????:                           f_lzc = 24;
            32'b1????????:                          f_lzc = 23;
            32'b1?????????:                         f_lzc = 22;
            32'b1??????????:                        f_lzc = 21;
            32'b1???????????:                       f_lzc = 20;
            32'b1????????????:                      f_lzc = 19;
            32'b1?????????????:                     f_lzc = 18;
            32'b1??????????????:                    f_lzc = 17;
            32'b1???????????????:                   f_lzc = 16;
            32'b1????????????????:                  f_lzc = 15;
            32'b1?????????????????:                 f_lzc = 14;
            32'b1??????????????????:                f_lzc = 13;
            32'b1???????????????????:               f_lzc = 12;
            32'b1????????????????????:              f_lzc = 11;
            32'b1?????????????????????:             f_lzc = 10;
            32'b1??????????????????????:            f_lzc = 9;
            32'b1???????????????????????:           f_lzc = 8;
            32'b1????????????????????????:          f_lzc = 7;
            32'b1?????????????????????????:         f_lzc = 6;
            32'b1??????????????????????????:        f_lzc = 5;
            32'b1???????????????????????????:       f_lzc = 4;
            32'b1????????????????????????????:      f_lzc = 3;
            32'b1?????????????????????????????:     f_lzc = 2;
            32'b1??????????????????????????????:    f_lzc = 1;
            default:                                f_lzc = 0;
        endcase
    endfunction

    assign lzc_cnt = f_lzc(i_data);

endmodule




//module lzc#(int WIDTH=8)
//  (input wire[WIDTH-1:0] i_data,
//   output wire [$clog2(WIDTH):0] lzc_cnt
//   );
//
//   wire       allzeroes;
//
//   function bit f(bit[WIDTH-1:0] x, int size);
//      bit                        jval = 0;
//      bit                        ival = 0;
//
//      for(int i = 1; i < size; i+=2) begin
//         jval = 1;
//         for(int j = i+1; j < size; j+=2) begin
//            jval &= ~x[j];
//         end
//         ival |= jval & x[i];
//      end
//
//      return ival;
//
//   endfunction // f
//
//   function bit[WIDTH-1:0] f_input(bit[WIDTH-1:0] x, int stage );
//      bit[WIDTH-1:0] dout = 0;
//      int            stagePow2 = 2**stage;
//      int            j=0;
//      for(int i=0; i<WIDTH; i++) begin
//         dout[j] |= x[i];
//         if(i % stagePow2 == stagePow2 - 1)
//           j++;
//      end
//      return dout;
//   endfunction
//
//   genvar i;
//
//   assign allzeroes = ~(|i_data);
//
//   assign lzc_cnt[$clog2(WIDTH)] = allzeroes;
//
//   generate
//      for(i=0; i < $clog2(WIDTH); i++) begin
//         assign lzc_cnt[i] = ~allzeroes & ~f(f_input(i_data, i),WIDTH);
//      end
//   endgenerate
//
//endmodule
